library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity BROM_TW is
    port(
        clk : in std_logic;
        raddr: in std_logic_vector(8 downto 0);
        dout: out std_logic_vector(15 downto 0)
    );
end entity BROM_TW;

architecture RTL of BROM_TW is
    -- brom
    type rom_type is array (0 to 256) of std_logic_vector(15 downto 0);
    signal rom: rom_type;
begin

    -- read operation
    process(clk)
    begin
        if rising_edge(clk) then
            case(raddr) is
                when "000000000" => dout <= x"fbec";
                when "000000001" => dout <= x"fd0a";
                when "000000010" => dout <= x"fe99";
                when "000000011" => dout <= x"fa13";
                when "000000100" => dout <= x"05d5";
                when "000000101" => dout <= x"058e";
                when "000000110" => dout <= x"011f";
                when "000000111" => dout <= x"00ca";
                when "000001000" => dout <= x"ff55";
                when "000001001" => dout <= x"026e";
                when "000001010" => dout <= x"0629";
                when "000001011" => dout <= x"00b6";
                when "000001100" => dout <= x"03c2";
                when "000001101" => dout <= x"fb4e";
                when "000001110" => dout <= x"fa3e";
                when "000001111" => dout <= x"05bc";
                when "000010000" => dout <= x"023d";
                when "000010001" => dout <= x"fad3";
                when "000010010" => dout <= x"0108";
                when "000010011" => dout <= x"017f";
                when "000010100" => dout <= x"fcc3";
                when "000010101" => dout <= x"05b2";
                when "000010110" => dout <= x"f9be";
                when "000010111" => dout <= x"ff7e";
                when "000011000" => dout <= x"fd57";
                when "000011001" => dout <= x"03f9";
                when "000011010" => dout <= x"02dc";
                when "000011011" => dout <= x"0260";
                when "000011100" => dout <= x"f9fa";
                when "000011101" => dout <= x"019b";
                when "000011110" => dout <= x"ff33";
                when "000011111" => dout <= x"f9dd";
                when "000100000" => dout <= x"04c7";
                when "000100001" => dout <= x"028c";
                when "000100010" => dout <= x"fdd8";
                when "000100011" => dout <= x"03f7";
                when "000100100" => dout <= x"faf3";
                when "000100101" => dout <= x"05d3";
                when "000100110" => dout <= x"fee6";
                when "000100111" => dout <= x"f9f8";
                when "000101000" => dout <= x"0204";
                when "000101001" => dout <= x"fff8";
                when "000101010" => dout <= x"fec0";
                when "000101011" => dout <= x"fd66";
                when "000101100" => dout <= x"f9ae";
                when "000101101" => dout <= x"fb76";
                when "000101110" => dout <= x"007e";
                when "000101111" => dout <= x"05bd";
                when "000110000" => dout <= x"fcab";
                when "000110001" => dout <= x"ffa6";
                when "000110010" => dout <= x"fef1";
                when "000110011" => dout <= x"033e";
                when "000110100" => dout <= x"006b";
                when "000110101" => dout <= x"fa73";
                when "000110110" => dout <= x"ff09";
                when "000110111" => dout <= x"fc49";
                when "000111000" => dout <= x"fe72";
                when "000111001" => dout <= x"03c1";
                when "000111010" => dout <= x"fa1c";
                when "000111011" => dout <= x"fd2b";
                when "000111100" => dout <= x"01c0";
                when "000111101" => dout <= x"fbd7";
                when "000111110" => dout <= x"02a5";
                when "000111111" => dout <= x"fb05";
                when "001000000" => dout <= x"fbb1";
                when "001000001" => dout <= x"01ae";
                when "001000010" => dout <= x"022b";
                when "001000011" => dout <= x"034b";
                when "001000100" => dout <= x"fb1d";
                when "001000101" => dout <= x"0367";
                when "001000110" => dout <= x"060e";
                when "001000111" => dout <= x"0069";
                when "001001000" => dout <= x"01a6";
                when "001001001" => dout <= x"024b";
                when "001001010" => dout <= x"00b1";
                when "001001011" => dout <= x"ff15";
                when "001001100" => dout <= x"fedd";
                when "001001101" => dout <= x"fe34";
                when "001001110" => dout <= x"0626";
                when "001001111" => dout <= x"0675";
                when "001010000" => dout <= x"ff0a";
                when "001010001" => dout <= x"030a";
                when "001010010" => dout <= x"0487";
                when "001010011" => dout <= x"ff6d";
                when "001010100" => dout <= x"fcf7";
                when "001010101" => dout <= x"05cb";
                when "001010110" => dout <= x"fda6";
                when "001010111" => dout <= x"045f";
                when "001011000" => dout <= x"f9ca";
                when "001011001" => dout <= x"0284";
                when "001011010" => dout <= x"fc98";
                when "001011011" => dout <= x"015d";
                when "001011100" => dout <= x"01a2";
                when "001011101" => dout <= x"0149";
                when "001011110" => dout <= x"ff64";
                when "001011111" => dout <= x"ffb5";
                when "001100000" => dout <= x"0331";
                when "001100001" => dout <= x"0449";
                when "001100010" => dout <= x"025b";
                when "001100011" => dout <= x"0262";
                when "001100100" => dout <= x"052a";
                when "001100101" => dout <= x"fafb";
                when "001100110" => dout <= x"fa47";
                when "001100111" => dout <= x"0180";
                when "001101000" => dout <= x"fb41";
                when "001101001" => dout <= x"ff78";
                when "001101010" => dout <= x"04c2";
                when "001101011" => dout <= x"fac9";
                when "001101100" => dout <= x"fc96";
                when "001101101" => dout <= x"00dc";
                when "001101110" => dout <= x"fb5d";
                when "001101111" => dout <= x"f985";
                when "001110000" => dout <= x"fb5f";
                when "001110001" => dout <= x"fa06";
                when "001110010" => dout <= x"fb02";
                when "001110011" => dout <= x"031a";
                when "001110100" => dout <= x"fa1a";
                when "001110101" => dout <= x"fcaa";
                when "001110110" => dout <= x"fc9a";
                when "001110111" => dout <= x"01de";
                when "001111000" => dout <= x"ff94";
                when "001111001" => dout <= x"fecc";
                when "001111010" => dout <= x"03e4";
                when "001111011" => dout <= x"03df";
                when "001111100" => dout <= x"03be";
                when "001111101" => dout <= x"fa4c";
                when "001111110" => dout <= x"05f2";
                when "001111111" => dout <= x"065c";
                ----------------------------------
                when "010000010" => dout <= x"FBB1";
                when "010000011" => dout <= x"044F";
                when "010000100" => dout <= x"01AE";
                when "010000101" => dout <= x"FE52";
                when "010000110" => dout <= x"022B";
                when "010000111" => dout <= x"FDD5";
                when "010001000" => dout <= x"034B";
                when "010001001" => dout <= x"FCB5";
                when "010001010" => dout <= x"FB1D";
                when "010001011" => dout <= x"04E3";
                when "010001100" => dout <= x"0367";
                when "010001101" => dout <= x"FC99";
                when "010001110" => dout <= x"060E";
                when "010001111" => dout <= x"F9F2";
                when "010010000" => dout <= x"0069";
                when "010010001" => dout <= x"FF97";
                when "010010010" => dout <= x"01A6";
                when "010010011" => dout <= x"FE5A";
                when "010010100" => dout <= x"024B";
                when "010010101" => dout <= x"FDB5";
                when "010010110" => dout <= x"00B1";
                when "010010111" => dout <= x"FF4F";
                when "010011000" => dout <= x"FF15";
                when "010011001" => dout <= x"00EB";
                when "010011010" => dout <= x"FEDD";
                when "010011011" => dout <= x"0123";
                when "010011100" => dout <= x"FE34";
                when "010011101" => dout <= x"01CC";
                when "010011110" => dout <= x"0626";
                when "010011111" => dout <= x"F9DA";
                when "010100000" => dout <= x"0675";
                when "010100001" => dout <= x"F98B";
                when "010100010" => dout <= x"FF0A";
                when "010100011" => dout <= x"00F6";
                when "010100100" => dout <= x"030A";
                when "010100101" => dout <= x"FCF6";
                when "010100110" => dout <= x"0487";
                when "010100111" => dout <= x"FB79";
                when "010101000" => dout <= x"FF6D";
                when "010101001" => dout <= x"0093";
                when "010101010" => dout <= x"FCF7";
                when "010101011" => dout <= x"0309";
                when "010101100" => dout <= x"05CB";
                when "010101101" => dout <= x"FA35";
                when "010101110" => dout <= x"FDA6";
                when "010101111" => dout <= x"025A";
                when "010110000" => dout <= x"045F";
                when "010110001" => dout <= x"FBA1";
                when "010110010" => dout <= x"F9CA";
                when "010110011" => dout <= x"0636";
                when "010110100" => dout <= x"0284";
                when "010110101" => dout <= x"FD7C";
                when "010110110" => dout <= x"FC98";
                when "010110111" => dout <= x"0368";
                when "010111000" => dout <= x"015D";
                when "010111001" => dout <= x"FEA3";
                when "010111010" => dout <= x"01A2";
                when "010111011" => dout <= x"FE5E";
                when "010111100" => dout <= x"0149";
                when "010111101" => dout <= x"FEB7";
                when "010111110" => dout <= x"FF64";
                when "010111111" => dout <= x"009C";
                when "011000000" => dout <= x"FFB5";
                when "011000001" => dout <= x"004B";
                when "011000010" => dout <= x"0331";
                when "011000011" => dout <= x"FCCF";
                when "011000100" => dout <= x"0449";
                when "011000101" => dout <= x"FBB7";
                when "011000110" => dout <= x"025B";
                when "011000111" => dout <= x"FDA5";
                when "011001000" => dout <= x"0262";
                when "011001001" => dout <= x"FD9E";
                when "011001010" => dout <= x"052A";
                when "011001011" => dout <= x"FAD6";
                when "011001100" => dout <= x"FAFB";
                when "011001101" => dout <= x"0505";
                when "011001110" => dout <= x"FA47";
                when "011001111" => dout <= x"05B9";
                when "011010000" => dout <= x"0180";
                when "011010001" => dout <= x"FE80";
                when "011010010" => dout <= x"FB41";
                when "011010011" => dout <= x"04BF";
                when "011010100" => dout <= x"FF78";
                when "011010101" => dout <= x"0088";
                when "011010110" => dout <= x"04C2";
                when "011010111" => dout <= x"FB3E";
                when "011011000" => dout <= x"FAC9";
                when "011011001" => dout <= x"0537";
                when "011011010" => dout <= x"FC96";
                when "011011011" => dout <= x"036A";
                when "011011100" => dout <= x"00DC";
                when "011011101" => dout <= x"FF24";
                when "011011110" => dout <= x"FB5D";
                when "011011111" => dout <= x"04A3";
                when "011100000" => dout <= x"F985";
                when "011100001" => dout <= x"067B";
                when "011100010" => dout <= x"FB5F";
                when "011100011" => dout <= x"04A1";
                when "011100100" => dout <= x"FA06";
                when "011100101" => dout <= x"05FA";
                when "011100110" => dout <= x"FB02";
                when "011100111" => dout <= x"04FE";
                when "011101000" => dout <= x"031A";
                when "011101001" => dout <= x"FCE6";
                when "011101010" => dout <= x"FA1A";
                when "011101011" => dout <= x"05E6";
                when "011101100" => dout <= x"FCAA";
                when "011101101" => dout <= x"0356";
                when "011101110" => dout <= x"FC9A";
                when "011101111" => dout <= x"0366";
                when "011110000" => dout <= x"01DE";
                when "011110001" => dout <= x"FE22";
                when "011110010" => dout <= x"FF94";
                when "011110011" => dout <= x"006C";
                when "011110100" => dout <= x"FECC";
                when "011110101" => dout <= x"0134";
                when "011110110" => dout <= x"03E4";
                when "011110111" => dout <= x"FC1C";
                when "011111000" => dout <= x"03DF";
                when "011111001" => dout <= x"FC21";
                when "011111010" => dout <= x"03BE";
                when "011111011" => dout <= x"FC42";
                when "011111100" => dout <= x"FA4C";
                when "011111101" => dout <= x"05B4";
                when "011111110" => dout <= x"05F2";
                when "011111111" => dout <= x"FA0E";
                when "100000000" => dout <= x"065C";
                when "100000001" => dout <= x"F9A4";    
                when others => dout <= x"0000";
            end case;
        end if;
    end process;
end architecture RTL;